*****************************************************************************************************************************************
*SRC=DMMT3906;DI_DMMT3906;BJTs PNP; Si;  40.0V  0.200A  257MHz   Diodes Inc. Matched BJTs - Single device of dual
.MODEL DI_DMMT3906  PNP (IS=20.3f NF=1.00 BF=437 VAF=114
+ IKF=44.6m ISE=6.81p NE=2.00 BR=4.00 NR=1.00
+ VAR=20.0 IKR=0.120 RE=1.16 RB=4.63 RC=0.463
+ XTB=1.5 CJE=23.5p VJE=1.10 MJE=0.500 CJC=10.7p VJC=0.300
+ MJC=0.300 TF=504p TR=94.3n EG=1.12 )
*****************************************************************************************************************************************